module and_gate(output out1, input in1, in2);

  and (out1, in1, in2);

endmodule

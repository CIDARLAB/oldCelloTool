module NOT(A,Y);
   input A;
   output Y;
endmodule // NOT
module NOR(A,B,Y);
   input A;
   input B;
   output Y;
endmodule // NOR
module DFF(C,D,Q);
   input C;
   input D;
   output Q;
endmodule // DFF
